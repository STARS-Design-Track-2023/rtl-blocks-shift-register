module shift_reg
#(
    parameter NUM_BITS = 8
) 
(
    input  logic                  clk, nrst, D,
    input  logic [1:0]            mode_i,
    input  logic [(NUM_BITS-1):0] par_i,
    output logic [(NUM_BITS-1):0] P
);

    // Write code here
    
endmodule
