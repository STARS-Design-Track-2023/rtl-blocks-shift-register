module shift_reg
(
    input  logic       clk, nrst, D,
    input  logic [1:0] mode_i,
    input  logic [7:0] par_i,
    output logic [7:0] P
);

    // Write code here
    
endmodule
